`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:49:25 10/03/2017 
// Design Name: 
// Module Name:    Floatingmul 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Floatingmul(
	output [31:0] out,
	input [31:0] A,
	input [31:0] B,
	input clk
    );
//mul m1();

endmodule
